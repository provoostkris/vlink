------------------------------------------------------------------------------
--  package for the nco designs
--  rev. 1.0 : 2025 Provoost Kris
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

package pckg_nco is

end pckg_nco;

package body pckg_nco is


end pckg_nco;