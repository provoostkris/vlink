------------------------------------------------------------------------------
--  package for the bpsk designs
--  rev. 1.0 : 2023 Provoost Kris
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

package pckg_bpsk_demod is


end pckg_bpsk_demod;

package body pckg_bpsk_demod is


end pckg_bpsk_demod;