------------------------------------------------------------------------------
--  package for the convolutional encoder
--  rev. 1.0 : 2023 Provoost Kris
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

package pckg_conv_enc is

end pckg_conv_enc;

package body pckg_conv_enc is
 
   
end pckg_conv_enc;