------------------------------------------------------------------------------
--  package for the bpsk_mod designs
--  rev. 1.0 : 2023 Provoost Kris
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

package pckg_bpsk_mod is


end pckg_bpsk_mod;

package body pckg_bpsk_mod is


end pckg_bpsk_mod;
