------------------------------------------------------------------------------
--  package for the pkt_asm functions
--  rev. 1.0 : 2025 Provoost Kris
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

package pckg_pkt_asm is


end pckg_pkt_asm;

package body pckg_pkt_asm is

end pckg_pkt_asm;