------------------------------------------------------------------------------
--  package for the bpsk designs
--  rev. 1.0 : 2023 Provoost Kris
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

package pckg_bpsk is


end pckg_bpsk;

package body pckg_bpsk is


end pckg_bpsk;
