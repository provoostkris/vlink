------------------------------------------------------------------------------
--  TOP level design file for virtual link
--  rev. 1.0 : 2022 Provoost Kris
------------------------------------------------------------------------------

library ieee;
use     ieee.std_logic_1164.all;
use     ieee.numeric_std.all;

entity vlink is
	generic(
	);
	port(
	);
end entity vlink;

architecture rtl of vlink is

begin

end architecture rtl;