------------------------------------------------------------------------------
--  package for the crc functions
--  rev. 1.0 : 2023 Provoost Kris
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

package pckg_dac is

end pckg_dac;

package body pckg_dac is


end pckg_dac;