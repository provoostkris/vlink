------------------------------------------------------------------------------
--  package for the sei designs
--  rev. 1.0 : 2022 Provoost Kris
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

package pckg_sei is


end pckg_sei;

package body pckg_sei is


end pckg_sei;